module adder(input logic[11:0] a,
             input logic [11:0] b,
             output logic[11:0] y);
                assign y= a+b;
endmodule